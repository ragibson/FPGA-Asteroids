`timescale 1ns / 1ps
`default_nettype none

module top #(
    //parameter imem_init="imem_screentest.mem",        // use this line for synthesis/board deployment
    parameter imem_init="imem_screentest_nopause.mem",  // use this line for simulation/testing
    parameter dmem_init="dmem_screentest.mem",          // file to initialize data memory
    parameter smem_init="smem_screentest.mem",          // file to initialize screen memory
    parameter bmem_init="bmem_screentest.mem"           // file to initialize bitmap memory
)(
    input wire clk, reset,
    input wire ps2_data,
    input wire ps2_clk,
    input wire aclMISO,
    output wire aclSCK,
    output wire aclMOSI,
    output wire aclSS,
    output wire audPWM,
    output wire audEn,
    output wire [15:0] LED,
    output wire [7:0] segments,
    output wire [7:0] digitselect,
    output wire [3:0] red, green, blue,
    output wire hsync, vsync
);
   wire [31:0] pc, instr, mem_readdata, mem_writedata, mem_addr;
   wire mem_wr;
   wire clk100, clk50, clk25, clk12;
   
   wire [10:0] smem_addr;
   wire [11:0] bmem_color;
   wire unsigned [31:0] period;
   wire [1:0] charcode;
   wire [31:0] keyb_char;
   wire enable = 1'b1;      // we will use this later for debugging
   assign audEn = 1'b1;

   // Uncomment *only* one of the following two lines:
   //    when synthesizing, use the first line
   //    when simulating, get rid of the clock divider, and use the second line
   //
   //clockdivider_Nexys4 clkdv(clk, clk100, clk50, clk25, clk12);   // use this line for synthesis/board deployment
   assign clk100=clk; assign clk50=clk; assign clk25=clk; assign clk12=clk;  // use this line for simulation/testing

   // For synthesis:  use an appropriate clock frequency(ies) below
   //   clk100 will work for hardly anyone
   //   clk50 or clk 25 may work for some
   //   clk12 should work for everyone!  So, please use clk12 for your processor and data memory.
   //
   // Important:  Use the same clock frequency for the MIPS and the memIO modules.
   // The I/O devices, however, should keep the 100 MHz clock.
   // For example:

   mips mips(clk12, reset, enable, pc, instr, mem_wr, mem_addr, mem_writedata, mem_readdata);
   rom_module #(.Nloc(256), .Dbits(32), .initfile(imem_init)) imem(pc[31:2], instr);
   memIO #(.Nloc(64), .Dbits(32), .numChars(4), .dmem_init(dmem_init), .smem_init(smem_init)) memIO
          (clk12, mem_wr, mem_addr, mem_writedata, smem_addr, accelX, accelY, keyb_char, mem_readdata, LED, period, charcode);

   // I/O devices
   //
   // Note: All I/O devices were developed assuming a 100 MHz clock.
   //   Therefore, the clock sent to them must be clk100, not any of the
   //   slower clocks generated by the clock divider.

   vgadisplaydriver #(.numChars(4), .initfile(bmem_init)) display
                     (clk100, charcode, smem_addr, bmem_color, red, green, blue, hsync, vsync);

   // Uncomment the following to instantiate these other I/O devices.
   //   You will have to declare all the wires that connect to them.
   //
   wire [8:0] accelX, accelY;
   wire [11:0] accelTmp;
   keyboard keyb(clk100, ps2_clk, ps2_data, keyb_char);
   display8digit disp(keyb_char, clk100, segments, digitselect);
   accelerometer accel(clk100, aclSCK, aclMOSI, aclMISO, aclSS, accelX, accelY, accelTmp);
   montek_sound_Nexys4 sound(clk100, period, audPWM);

endmodule

